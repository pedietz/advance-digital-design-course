
module diffeq (
    output signed y[8:0];
    input  signed x[8:0];
);
    
endmodule